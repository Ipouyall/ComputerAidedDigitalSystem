`timescale 1ns/1ns
module  LUT(clk, addr, q);
    input [4:0] addr ;
    input clk;
    output reg [63:0] q; 
    always@(posedge clk) begin 
        case(addr) 
            0: q <= 64'h0000000000000001;
            1: q <= 64'h0000000000008082;
            2: q <= 64'h800000000000808a;
            3: q <= 64'h8000000080008000;
            4: q <= 64'h000000000000808b;
            5: q <= 64'h0000000080000001;
            6: q <= 64'h8000000080008081;
            7: q <= 64'h8000000000008009;
            8: q <= 64'h000000000000008a;
            9: q <= 64'h0000000000000088;
            10:q <= 64'h0000000080008009;
            11:q <= 64'h000000008000000a;
            12: q <= 64'h000000008000808b;
            13: q <= 64'h800000000000008b;
            14: q <= 64'h8000000000008089;
            15: q <= 64'h8000000000008003;
            16: q <= 64'h8000000000008002;
            17: q <= 64'h8000000000000080;
            18: q <= 64'h000000000000800a;
            19: q <= 64'h800000008000000a;
            20: q <= 64'h8000000080008081;
            21: q <= 64'h8000000000008080;
            22: q <= 64'h0000000080000001;
            23: q <= 64'h8000000080008008;
            default:q <= 64'h00;
        endcase 
    end
endmodule


